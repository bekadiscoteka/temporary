Vim�UnDo� qE=uO;֨����_�������5n���#%�   �   `include "top_assist/bin2bcd.v"            ;       ;   ;   ;    h:�    _�                     *        ����                                                                                                                                                                                                                                                                                                                            w          *           v        h�F     �   )   +   �   N   +	always @(posedge clk, posedge reset) begin   		if (reset) begin   		   enable <= 4'b0000;	   			state <= 0;   			start <= 0;   		end   		case (state)    			IDLE: begin   				start <= 0;   				if (read) begin   					enable <= 4'b0100;   					state <= PROC;	   				end   			end   			PROC: begin   				if (read) begin   !					if (enable == 4'b0001) begin   						if (ascii != 45) begin   							enable <= 0;   							start <= 1;   							state <= IDLE;   							end   					end   					else begin   3						enable <= ascii == 45 ? enable : enable >> 1;   					end   				end   			end	   			endcase   	end	       +	always @(posedge clk, posedge reset) begin   		if (reset) begin   
			a <= 0;   
			b <= 0;   
			c <= 0;   
			d <= 0;   			temp <= 0;   		end   		else if (read) begin   			if (enable[2]) begin   				if (ascii == 45) begin   				   	temp <= 1;   				end   				else begin   ,					b <= temp ? -(ascii - 48) : ascii - 48;   					temp <= 0;   				end	   			end   			else if (enable[1]) begin   				if (ascii == 45) begin   				   	temp <= 1;   				end   				else begin   ,					c <= temp ? -(ascii - 48) : ascii - 48;   					temp <= 0;   				end	   			end   			else if (enable[0]) begin   				if (ascii == 45) begin   				   	temp <= 1;   				end   				else begin   ,					d <= temp ? -(ascii - 48) : ascii - 48;   					temp <= 0;   				end	   			end   			else begin   				if (ascii == 45) begin   				   	temp <= 1;   				end   				else begin   ,					a <= temp ? -(ascii - 48) : ascii - 48;   					temp <= 0;   				end   			end   		end   	end5�_�                    *        ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�G     �   )   ,   p       5�_�                    *       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�Q     �   *   -   r      		�   *   ,   q    5�_�                    +       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�^     �   +   .   t      			�   +   -   s    5�_�                    ,   	    ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�s     �   ,   /   v      				�   ,   .   u    5�_�                    -       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�z     �   -   /   x      					�   -   /   w    5�_�                    .   	    ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   -   /   x      						if (5�_�      	              .       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   -   5   x      					�   .   /   x    5�_�      
           	   /       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   .   0   ~      				   	temp <= 1;5�_�   	              
   0       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   /   1   ~      				end5�_�   
                 1       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   0   2   ~      				else begin5�_�                    2       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   1   3   ~      ,					b <= temp ? -(ascii - 48) : ascii - 48;5�_�                    3       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   2   4   ~      					temp <= 0;5�_�                    4       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�    �   3   5   ~      				end5�_�                    2       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h��     �   1   3   ~      -						b <= temp ? -(ascii - 48) : ascii - 48;5�_�                    2       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h��     �   1   3   ~      -						1 <= temp ? -(ascii - 48) : ascii - 48;5�_�                    3       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h��     �   3   5         						�   3   5   ~    5�_�                    6       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h��     �   6   9   �      				�   6   8       5�_�                    7       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h��     �   7   9   �      					�   7   9   �    5�_�                    8       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h��     �   7   ?   �      						�   8   9   �    5�_�                    9       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h��     �   8   :   �      				   	temp <= 1;5�_�                    :       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�      �   9   ;   �      				end5�_�                    ;       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   :   <   �      				else begin5�_�                    <       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   ;   =   �      ,					b <= temp ? -(ascii - 48) : ascii - 48;5�_�                    =       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   <   >   �      					temp <= 0;5�_�                    >       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�    �   =   ?   �      				end	5�_�                    =       ����                                                                                                                                                                                                                                                                                                                            *          *           v        h�     �   =   ?   �      						�   =   ?   �    5�_�                    @        ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�     �   @   C   �      				�   @   B   �    5�_�                    A       ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�%     �   A   C   �    5�_�      !              A        ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�*     �   A   C   �      					�   A   C   �    5�_�      "           !   C        ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�9     �   B   K   �       �   C   D   �    5�_�   !   #           "   B        ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�>     �   A   B          						5�_�   "   $           #   F       ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�C     �   E   G   �      -						b <= temp ? -(ascii - 48) : ascii - 48;5�_�   #   %           $   H       ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�E     �   G   I   �      						state <= SET_C;5�_�   $   &           %   H       ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�G    �   G   I   �      						state <= SET_c;5�_�   %   '           &   J        ����                                                                                                                                                                                                                                                                                                                            I          B           v        h�N     �   J   M   �      				�   J   L   �    5�_�   &   (           '   K       ����                                                                                                                                                                                                                                                                                                                            I          B           v        h�T     �   K   M   �    5�_�   '   )           (   L        ����                                                                                                                                                                                                                                                                                                                            I          B           v        h�Z     �   K   T   �       �   L   M   �    5�_�   (   *           )   P       ����                                                                                                                                                                                                                                                                                                                            I          B           v        h�`    �   O   Q   �      -						c <= temp ? -(ascii - 48) : ascii - 48;5�_�   )   +           *   R       ����                                                                                                                                                                                                                                                                                                                            I          B           v        h�q     �   Q   S   �      						state <= SET_D;5�_�   *   ,           +   R       ����                                                                                                                                                                                                                                                                                                                            I          B           v        h�s    �   R   T   �      						�   R   T   �    5�_�   +   -           ,   -       ����                                                                                                                                                                                                                                                                                                                            I          B           v        h��   	 �   -   /   �      					�   -   /   �    5�_�   ,   .           -   X       ����                                                                                                                                                                                                                                                                                                                            J          C           v        h��   
 �   X   Z   �      		�   X   Z   �    5�_�   -   /           .   *       ����                                                                                                                                                                                                                                                                                                                            J          C           v        h��     �   *   -   �      		�   *   ,   �    5�_�   .   0           /   +       ����                                                                                                                                                                                                                                                                                                                            L          E           v        h��     �   +   /   �      			�   +   -   �    5�_�   /   1           0   %       ����                                                                                                                                                                                                                                                                                                                            O          H           v        h�    �   $   %          	reg [3:0] enable;5�_�   0   2           1   -       ����                                                                                                                                                                                                                                                                                                                            N          G           v        h�    �   -   2   �      			�   -   /   �    5�_�   1   3           2   %       ����                                                                                                                                                                                                                                                                                                                            R          K           v        h�    �   $   &   �      	reg state;5�_�   2   4           3          ����                                                                                                                                                                                                                                                                                                                            R          K           v        h�?     �                	parameter	IDLE=0,5�_�   3   5           4          ����                                                                                                                                                                                                                                                                                                                            Q          J           v        h�@     �                					PROC=1;5�_�   4   6           5          ����                                                                                                                                                                                                                                                                                                                            P          I           v        h�B    �         �      			5�_�   5   7           6          ����                                                                                                                                                                                                                                                                                                                            S          L           v        h�_    �         �    5�_�   6   8           7      
    ����                                                                                                                                                                                                                                                                                                                                                             h9�     �         �       `include "bcd2sseg_active_low.v"5�_�   7   9           8      
    ����                                                                                                                                                                                                                                                                                                                                                             h9�    �         �      `include "bin2bcd.v"5�_�   8   :           9          ����                                                                                                                                                                                                                                                                                                                                                             h:�     �         �      +`include "top_assist/bcd2sseg_active_low.v"5�_�   9   ;           :          ����                                                                                                                                                                                                                                                                                                                                                             h:�     �         �      `include "top_assist/bin2bcd.v"5�_�   :               ;          ����                                                                                                                                                                                                                                                                                                                                                             h:�    �         �       `include "top_support/bin2bcd.v"5�_�             !       B        ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�4     �   B   C   �    �   A   C   �      						if (ascii == 45) begin   				   		temp <= 1;   					end   					else begin   -						b <= temp ? -(ascii - 48) : ascii - 48;   						temp <= 0;   						state <= SET_C;   					end						5�_�                     B       ����                                                                                                                                                                                                                                                                                                                            ?          8           v        h�0     �   B   C   �    �   A   C   �       										if (ascii == 45) begin   				   		temp <= 1;   					end   					else begin   -						b <= temp ? -(ascii - 48) : ascii - 48;   						temp <= 0;   						state <= SET_C;   
					end		5��