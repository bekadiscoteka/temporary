Vim�UnDo� ����ǋ���~
�k �5Z�}�/ޞ����   g   :	always @(posedge top.read) $display("read 1: %d", $time);   (   0      +       +   +   +    hc�   ) _�                     +       ����                                                                                                                                                                                                                                                                                                                            2          +          v       hUk     �   *   ,   l      F	always @(posedge top.divided_clk_tick) $display("%d %d %d %d %d %d ",   		top.bcd_set[(6*4)-1:(5*4)],   		top.bcd_set[(5*4)-1:(4*4)],   		top.bcd_set[(4*4)-1:(3*4)],   		top.bcd_set[(3*4)-1:(2*4)],   		top.bcd_set[(2*4)-1:(1*4)],   		top.bcd_set[(1*4)-1:(0*4)]   	);5�_�                    +       ����                                                                                                                                                                                                                                                                                                                            +          +          v       hUl     �   *   +          	always @(posedge5�_�                    *        ����                                                                                                                                                                                                                                                                                                                            +          +          v       hUl     �   )   *           5�_�                    *        ����                                                                                                                                                                                                                                                                                                                            *          *          v       hUm    �   )   *           5�_�                    %       ����                                                                                                                                                                                                                                                                                                                            *          *          v       hU~    �   $   %          		.banner_write(being_written)5�_�      
              $   !    ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�    �   #   %   a      !		.baund_rate_ready(baund_ready),5�_�                
   7       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�   	 �   6   8   a      		terminal="w";5�_�   
                 B       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�   
 �   A   C   a      		terminal="4";5�_�                    G       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�    �   F   H   a      		terminal="0";5�_�                    J       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�     �   J   L   b      		�   J   L   a    5�_�                    _       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�    �   ^   `   b      	   	5�_�                    _       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�    �   _   a   c      		�   _   a   b    5�_�                    _       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hVC     �   _   a   d      		�   _   a   c    5�_�                    `       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hV�    �   _   a   d      		wait(5�_�                    7       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h[�     �   6   8   d      		terminal="3";5�_�                    =       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h[�     �   <   >   d      		terminal="3";5�_�                    G       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h[�    �   F   H   d      		terminal="3";5�_�                    K       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h\[     �   J   K          		/*5�_�                    N       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h\k    �   N   P   d      		�   N   P   c    5�_�                    a       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h]    �   `   a          		#1000;5�_�                    a       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h]     �   `   b   c      		#30 $finish;	5�_�                    `       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h]%     �   `   c   d      		�   `   b   c    5�_�                    a        ����                                                                                                                                                                                                                                                                                                                            )          )          v       h]�     �   `   b   e       		$display("math expr is done");5�_�                    a       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h]�     �   `   b   e       		$display("math expr is done");5�_�                    b       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h]�    �   a   c   e      		wait(top.5�_�                    b       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h]�    �   b   d   f      		�   b   d   e    5�_�                    =       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h`�     �   <   >   f      		terminal="2";5�_�                     G       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h`�    �   F   H   f      		terminal="4";5�_�      !               b       ����                                                                                                                                                                                                                                                                                                                            )          )          v       h`�    �   b   d   g      		�   b   d   f    5�_�       "           !   c       ����                                                                                                                                                                                                                                                                                                                            )          )          v       ha     �   b   c          		#10;5�_�   !   #           "   c       ����                                                                                                                                                                                                                                                                                                                            )          )          v       ha    �   c   e   g      		�   c   e   f    5�_�   "   $           #   G       ����                                                                                                                                                                                                                                                                                                                            )          )          v       ha�    �   F   H   g      		terminal="-3";5�_�   #   %           $   G       ����                                                                                                                                                                                                                                                                                                                            )          )          v       ha�    �   F   H   g      		terminal="3";5�_�   $   &           %   O       ����                                                                                                                                                                                                                                                                                                                            )          )          v       ha�     �   N   O          		/*5�_�   %   '           &   Q       ����                                                                                                                                                                                                                                                                                                                            )          )          v       ha�    �   P   R   f      		terminal="4";5�_�   &   (           '   S   	    ����                                                                                                                                                                                                                                                                                                                            )          )          v       ha�   % �   S   U   g      		�   S   U   f    5�_�   '   )           (   '        ����                                                                                                                                                                                                                                                                                                                            )          )          v       hc�     �   '   *   h      	�   '   )   g    5�_�   (   *           )   )       ����                                                                                                                                                                                                                                                                                                                            +          +          v       hc�     �   (   )          	end5�_�   )   +           *   )        ����                                                                                                                                                                                                                                                                                                                            *          *          v       hc�   & �   '   )   h      !	always @(posedge top.read) begin    �   (   *   h       5�_�   *               +   (   0    ����                                                                                                                                                                                                                                                                                                                            )          )          v       hc�   ) �   '   )   g      :	always @(posedge top.read) $display("read 1: %d", $time);5�_�             
      7       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�    �   6   8   a      		terminal="3";5�_�      	              :   	    ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�    �   9   <        5�_�                  	   :       ����                                                                                                                                                                                                                                                                                                                            )          )          v       hU�    �   9   ;        5��