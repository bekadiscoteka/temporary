Vim�UnDo� �IJ-f�ʅ0�"�F6�V_��$͎���"*�,��   c                                  h{�    _�                     (       ����                                                                                                                                                                                                                                                                                                                                                             hy    �   (   *   h      	�   (   *   g    5�_�                    )       ����                                                                                                                                                                                                                                                                                                                                                             hyD    �   (   *   h      +	always @(posedge start) $display("start");5�_�                    7       ����                                                                                                                                                                                                                                                                                                                            ;   	       7          v       h{�     �   6   8   h      		#1;   		terminal="1";   
		write=1;   		@(posedge clk);   
		write=0;5�_�                     7       ����                                                                                                                                                                                                                                                                                                                            7          7          v       h{�    �   6   7          		5��